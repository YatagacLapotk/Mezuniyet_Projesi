`include "SABIT_VERILER/sabit_veriler.vh"
module MDU (
    input 
);
    
endmodule