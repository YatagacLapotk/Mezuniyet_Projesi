`ifndef sabit_veriler_VH
`define sabit_veriler_VH

`define ADDRESS_WIDTH 5
`define DATA_WIDTH 32
`define REG_FILE_DEPTH 32
`define INSTRUCTION_WIDTH 32
`define MUL_WIDTH 64
`define OPCODE_WIDTH 7
`define FUNCT3_WIDTH 3
`define FUNCT7_WIDTH 7




// MUL/DIV Operations
`define MUL    32'b0000001??????????000?????0110011
`define MULH   32'b0000001??????????001?????0110011
`define MULHU  32'b0000001??????????010?????0110011
`define MULHSU 32'b0000001??????????011?????0110011
`define DIV    32'b0000001??????????100?????0110011
`define DIVU   32'b0000001??????????101?????0110011
`define REM    32'b0000001??????????110?????0110011
`define REMU   32'b0000001??????????111?????0110011

`endif // sabit_veriler_VH

// RV32I Operations
`define LUI 32'b?????????????????????????0110111
`define AUIPC 32'b?????????????????????????0010111
`define JAL 32'b?????????????????????????1101111
`define JALR 32'b?????????????????000?????1100111
`define BEQ 32'b?????????????????000?????1100011
`define BNE 32'b?????????????????001?????1100011
`define BLT 32'b?????????????????100?????1100011
`define BGE 32'b?????????????????101?????1100011
`define BLTU 32'b?????????????????110?????1100011
`define BGEU 32'b?????????????????111?????1100011
`define LB 32'b?????????????????000?????0000011
`define LH 32'b?????????????????001?????0000011
`define LW 32'b?????????????????010?????0000011
`define LBU 32'b?????????????????100?????0000011
`define LHU 32'b?????????????????101?????0000011
`define SB 32'b?????????????????000?????0100011
`define SH 32'b?????????????????001?????0100011
`define SW 32'b?????????????????010?????0100011
`define ADDI 32'b?????????????????000?????0010011
`define SLTI 32'b?????????????????010?????0010011
`define SLTIU 32'b?????????????????011?????0010011
`define XORI 32'b?????????????????100?????0010011
`define ORI 32'b?????????????????110?????0010011
`define ANDI 32'b?????????????????111?????0010011
`define SLLI 32'b0000000??????????001?????0010011
`define SRLI 32'b0000000??????????101?????0010011
`define SRAI 32'b0100000??????????101?????0010011
`define ADD 32'b0000000??????????000?????0110011
`define SUB 32'b0100000??????????000?????0110011
`define SLL 32'b0000000??????????001?????0110011
`define SLT 32'b0000000??????????010?????0110011
`define SLTU 32'b0000000??????????011?????0110011
`define XOR 32'b0000000??????????100?????0110011
`define SRL 32'b0000000??????????101?????0110011
`define SRA 32'b0100000??????????101?????0110011
`define OR 32'b0000000??????????110?????0110011
`define AND 32'b0000000??????????111?????0110011