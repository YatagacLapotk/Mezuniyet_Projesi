module  (
    ports
);
    
endmodule