module REG_FILE_TB ();

wire          clk;
wire          res;
wire [4:0]    A1;
wire [4:0]    A2;
wire [4:0]    A3;
wire [31:0]   WD;
reg  [31:0]   RD1;
reg  [31:0]   RD2;

    
endmodule